// system_0.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module system_0 (
		output wire        audio_0_avalon_slave_0_export_oAUD_DATA,                     //           audio_0_avalon_slave_0_export.oAUD_DATA
		output wire        audio_0_avalon_slave_0_export_oAUD_LRCK,                     //                                        .oAUD_LRCK
		output wire        audio_0_avalon_slave_0_export_oAUD_BCK,                      //                                        .oAUD_BCK
		output wire        audio_0_avalon_slave_0_export_oAUD_XCK,                      //                                        .oAUD_XCK
		input  wire        audio_0_avalon_slave_0_export_iCLK_18_4,                     //                                        .iCLK_18_4
		input  wire [3:0]  button_pio_external_connection_export,                       //          button_pio_external_connection.export
		input  wire        clk_clk_in_clk,                                              //                              clk_clk_in.clk
		input  wire        clk_clk_in_reset_reset_n,                                    //                        clk_clk_in_reset.reset_n
		output wire [7:0]  led_green_external_connection_export,                        //           led_green_external_connection.export
		output wire [9:0]  led_red_external_connection_export,                          //             led_red_external_connection.export
		output wire        sd_clk_external_connection_export,                           //              sd_clk_external_connection.export
		inout  wire        sd_cmd_external_connection_export,                           //              sd_cmd_external_connection.export
		inout  wire        sd_dat_external_connection_export,                           //              sd_dat_external_connection.export
		output wire [11:0] sdram_0_wire_addr,                                           //                            sdram_0_wire.addr
		output wire [1:0]  sdram_0_wire_ba,                                             //                                        .ba
		output wire        sdram_0_wire_cas_n,                                          //                                        .cas_n
		output wire        sdram_0_wire_cke,                                            //                                        .cke
		output wire        sdram_0_wire_cs_n,                                           //                                        .cs_n
		inout  wire [15:0] sdram_0_wire_dq,                                             //                                        .dq
		output wire [1:0]  sdram_0_wire_dqm,                                            //                                        .dqm
		output wire        sdram_0_wire_ras_n,                                          //                                        .ras_n
		output wire        sdram_0_wire_we_n,                                           //                                        .we_n
		output wire [6:0]  seg7_display_conduit_end_oSEG0,                              //                seg7_display_conduit_end.oSEG0
		output wire [6:0]  seg7_display_conduit_end_oSEG1,                              //                                        .oSEG1
		output wire [6:0]  seg7_display_conduit_end_oSEG2,                              //                                        .oSEG2
		output wire [6:0]  seg7_display_conduit_end_oSEG3,                              //                                        .oSEG3
		output wire [6:0]  seg7_display_conduit_end_oSEG4,                              //                                        .oSEG4
		output wire [6:0]  seg7_display_conduit_end_oSEG5,                              //                                        .oSEG5
		output wire [6:0]  seg7_display_conduit_end_oSEG6,                              //                                        .oSEG6
		output wire [6:0]  seg7_display_conduit_end_oSEG7,                              //                                        .oSEG7
		inout  wire [15:0] sram_16bit_512k_0_avalon_slave_0_export_DQ,                  // sram_16bit_512k_0_avalon_slave_0_export.DQ
		output wire [17:0] sram_16bit_512k_0_avalon_slave_0_export_ADDR,                //                                        .ADDR
		output wire        sram_16bit_512k_0_avalon_slave_0_export_UB_N,                //                                        .UB_N
		output wire        sram_16bit_512k_0_avalon_slave_0_export_LB_N,                //                                        .LB_N
		output wire        sram_16bit_512k_0_avalon_slave_0_export_WE_N,                //                                        .WE_N
		output wire        sram_16bit_512k_0_avalon_slave_0_export_CE_N,                //                                        .CE_N
		output wire        sram_16bit_512k_0_avalon_slave_0_export_OE_N,                //                                        .OE_N
		input  wire [17:0] switch_pio_external_connection_export,                       //          switch_pio_external_connection.export
		inout  wire [7:0]  tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_data,     //         tri_state_bridge_0_bridge_0_out.tri_state_bridge_0_data
		output wire [0:0]  tri_state_bridge_0_bridge_0_out_write_n_to_the_cfi_flash_0,  //                                        .write_n_to_the_cfi_flash_0
		output wire [0:0]  tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_readn,    //                                        .tri_state_bridge_0_readn
		output wire [21:0] tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_address,  //                                        .tri_state_bridge_0_address
		output wire [0:0]  tri_state_bridge_0_bridge_0_out_select_n_to_the_cfi_flash_0, //                                        .select_n_to_the_cfi_flash_0
		input  wire        uart_0_external_connection_rxd,                              //              uart_0_external_connection.rxd
		output wire        uart_0_external_connection_txd                               //                                        .txd
	);

	wire         tri_state_bridge_0_pinsharer_0_tcm_request;                         // tri_state_bridge_0_pinSharer_0:request -> tri_state_bridge_0_bridge_0:request
	wire   [0:0] tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out; // tri_state_bridge_0_pinSharer_0:select_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0:tcs_select_n_to_the_cfi_flash_0
	wire  [21:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out;  // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_address -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_address
	wire   [0:0] tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out;  // tri_state_bridge_0_pinSharer_0:write_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0:tcs_write_n_to_the_cfi_flash_0
	wire         tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen;   // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data_outen -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data_outen
	wire   [7:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out;     // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data
	wire         tri_state_bridge_0_pinsharer_0_tcm_grant;                           // tri_state_bridge_0_bridge_0:grant -> tri_state_bridge_0_pinSharer_0:grant
	wire   [7:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in;      // tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data_in -> tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data_in
	wire   [0:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out;    // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_readn -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_readn
	wire         cfi_flash_0_tcm_data_outen;                                         // cfi_flash_0:tcm_data_outen -> tri_state_bridge_0_pinSharer_0:tcs0_data_outen
	wire         cfi_flash_0_tcm_request;                                            // cfi_flash_0:tcm_request -> tri_state_bridge_0_pinSharer_0:tcs0_request
	wire         cfi_flash_0_tcm_write_n_out;                                        // cfi_flash_0:tcm_write_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_write_n_out
	wire         cfi_flash_0_tcm_read_n_out;                                         // cfi_flash_0:tcm_read_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_read_n_out
	wire         cfi_flash_0_tcm_grant;                                              // tri_state_bridge_0_pinSharer_0:tcs0_grant -> cfi_flash_0:tcm_grant
	wire         cfi_flash_0_tcm_chipselect_n_out;                                   // cfi_flash_0:tcm_chipselect_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_chipselect_n_out
	wire  [21:0] cfi_flash_0_tcm_address_out;                                        // cfi_flash_0:tcm_address_out -> tri_state_bridge_0_pinSharer_0:tcs0_address_out
	wire   [7:0] cfi_flash_0_tcm_data_out;                                           // cfi_flash_0:tcm_data_out -> tri_state_bridge_0_pinSharer_0:tcs0_data_out
	wire   [7:0] cfi_flash_0_tcm_data_in;                                            // tri_state_bridge_0_pinSharer_0:tcs0_data_in -> cfi_flash_0:tcm_data_in
	wire  [31:0] nios2_qsys_0_data_master_readdata;                                  // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                               // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                               // nios2_qsys_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [24:0] nios2_qsys_0_data_master_address;                                   // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                      // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_readdatavalid;                             // mm_interconnect_0:nios2_qsys_0_data_master_readdatavalid -> nios2_qsys_0:d_readdatavalid
	wire         nios2_qsys_0_data_master_write;                                     // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                 // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                           // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                        // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [24:0] nios2_qsys_0_instruction_master_address;                            // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                               // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         nios2_qsys_0_instruction_master_readdatavalid;                      // mm_interconnect_0:nios2_qsys_0_instruction_master_readdatavalid -> nios2_qsys_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;           // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;        // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;            // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;               // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;              // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_seg7_display_avalon_slave_write;                  // mm_interconnect_0:SEG7_Display_avalon_slave_write -> SEG7_Display:iWR
	wire  [31:0] mm_interconnect_0_seg7_display_avalon_slave_writedata;              // mm_interconnect_0:SEG7_Display_avalon_slave_writedata -> SEG7_Display:iDIG
	wire         mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_chipselect;      // mm_interconnect_0:sram_16bit_512k_0_avalon_slave_0_chipselect -> sram_16bit_512k_0:iCE_N
	wire  [15:0] mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_readdata;        // sram_16bit_512k_0:oDATA -> mm_interconnect_0:sram_16bit_512k_0_avalon_slave_0_readdata
	wire  [17:0] mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_address;         // mm_interconnect_0:sram_16bit_512k_0_avalon_slave_0_address -> sram_16bit_512k_0:iADDR
	wire         mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_read;            // mm_interconnect_0:sram_16bit_512k_0_avalon_slave_0_read -> sram_16bit_512k_0:iOE_N
	wire   [1:0] mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_byteenable;      // mm_interconnect_0:sram_16bit_512k_0_avalon_slave_0_byteenable -> sram_16bit_512k_0:iBE_N
	wire         mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_write;           // mm_interconnect_0:sram_16bit_512k_0_avalon_slave_0_write -> sram_16bit_512k_0:iWE_N
	wire  [15:0] mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_writedata;       // mm_interconnect_0:sram_16bit_512k_0_avalon_slave_0_writedata -> sram_16bit_512k_0:iDATA
	wire  [15:0] mm_interconnect_0_audio_0_avalon_slave_0_readdata;                  // Audio_0:oDATA -> mm_interconnect_0:Audio_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_audio_0_avalon_slave_0_write;                     // mm_interconnect_0:Audio_0_avalon_slave_0_write -> Audio_0:iWR
	wire  [15:0] mm_interconnect_0_audio_0_avalon_slave_0_writedata;                 // mm_interconnect_0:Audio_0_avalon_slave_0_writedata -> Audio_0:iDATA
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata;            // nios2_qsys_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest;         // nios2_qsys_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess;         // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_debugaccess -> nios2_qsys_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address;             // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_address -> nios2_qsys_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read;                // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_read -> nios2_qsys_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable;          // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_byteenable -> nios2_qsys_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write;               // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_write -> nios2_qsys_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata;           // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_writedata -> nios2_qsys_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_epcs_controller_epcs_control_port_chipselect;     // mm_interconnect_0:epcs_controller_epcs_control_port_chipselect -> epcs_controller:chipselect
	wire  [31:0] mm_interconnect_0_epcs_controller_epcs_control_port_readdata;       // epcs_controller:readdata -> mm_interconnect_0:epcs_controller_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_controller_epcs_control_port_address;        // mm_interconnect_0:epcs_controller_epcs_control_port_address -> epcs_controller:address
	wire         mm_interconnect_0_epcs_controller_epcs_control_port_read;           // mm_interconnect_0:epcs_controller_epcs_control_port_read -> epcs_controller:read_n
	wire         mm_interconnect_0_epcs_controller_epcs_control_port_write;          // mm_interconnect_0:epcs_controller_epcs_control_port_write -> epcs_controller:write_n
	wire  [31:0] mm_interconnect_0_epcs_controller_epcs_control_port_writedata;      // mm_interconnect_0:epcs_controller_epcs_control_port_writedata -> epcs_controller:writedata
	wire         mm_interconnect_0_led_green_s1_chipselect;                          // mm_interconnect_0:led_green_s1_chipselect -> led_green:chipselect
	wire  [31:0] mm_interconnect_0_led_green_s1_readdata;                            // led_green:readdata -> mm_interconnect_0:led_green_s1_readdata
	wire   [1:0] mm_interconnect_0_led_green_s1_address;                             // mm_interconnect_0:led_green_s1_address -> led_green:address
	wire         mm_interconnect_0_led_green_s1_write;                               // mm_interconnect_0:led_green_s1_write -> led_green:write_n
	wire  [31:0] mm_interconnect_0_led_green_s1_writedata;                           // mm_interconnect_0:led_green_s1_writedata -> led_green:writedata
	wire         mm_interconnect_0_led_red_s1_chipselect;                            // mm_interconnect_0:led_red_s1_chipselect -> led_red:chipselect
	wire  [31:0] mm_interconnect_0_led_red_s1_readdata;                              // led_red:readdata -> mm_interconnect_0:led_red_s1_readdata
	wire   [1:0] mm_interconnect_0_led_red_s1_address;                               // mm_interconnect_0:led_red_s1_address -> led_red:address
	wire         mm_interconnect_0_led_red_s1_write;                                 // mm_interconnect_0:led_red_s1_write -> led_red:write_n
	wire  [31:0] mm_interconnect_0_led_red_s1_writedata;                             // mm_interconnect_0:led_red_s1_writedata -> led_red:writedata
	wire         mm_interconnect_0_sd_clk_s1_chipselect;                             // mm_interconnect_0:SD_CLK_s1_chipselect -> SD_CLK:chipselect
	wire  [31:0] mm_interconnect_0_sd_clk_s1_readdata;                               // SD_CLK:readdata -> mm_interconnect_0:SD_CLK_s1_readdata
	wire   [1:0] mm_interconnect_0_sd_clk_s1_address;                                // mm_interconnect_0:SD_CLK_s1_address -> SD_CLK:address
	wire         mm_interconnect_0_sd_clk_s1_write;                                  // mm_interconnect_0:SD_CLK_s1_write -> SD_CLK:write_n
	wire  [31:0] mm_interconnect_0_sd_clk_s1_writedata;                              // mm_interconnect_0:SD_CLK_s1_writedata -> SD_CLK:writedata
	wire         mm_interconnect_0_sd_cmd_s1_chipselect;                             // mm_interconnect_0:SD_CMD_s1_chipselect -> SD_CMD:chipselect
	wire  [31:0] mm_interconnect_0_sd_cmd_s1_readdata;                               // SD_CMD:readdata -> mm_interconnect_0:SD_CMD_s1_readdata
	wire   [1:0] mm_interconnect_0_sd_cmd_s1_address;                                // mm_interconnect_0:SD_CMD_s1_address -> SD_CMD:address
	wire         mm_interconnect_0_sd_cmd_s1_write;                                  // mm_interconnect_0:SD_CMD_s1_write -> SD_CMD:write_n
	wire  [31:0] mm_interconnect_0_sd_cmd_s1_writedata;                              // mm_interconnect_0:SD_CMD_s1_writedata -> SD_CMD:writedata
	wire         mm_interconnect_0_sd_dat_s1_chipselect;                             // mm_interconnect_0:SD_DAT_s1_chipselect -> SD_DAT:chipselect
	wire  [31:0] mm_interconnect_0_sd_dat_s1_readdata;                               // SD_DAT:readdata -> mm_interconnect_0:SD_DAT_s1_readdata
	wire   [1:0] mm_interconnect_0_sd_dat_s1_address;                                // mm_interconnect_0:SD_DAT_s1_address -> SD_DAT:address
	wire         mm_interconnect_0_sd_dat_s1_write;                                  // mm_interconnect_0:SD_DAT_s1_write -> SD_DAT:write_n
	wire  [31:0] mm_interconnect_0_sd_dat_s1_writedata;                              // mm_interconnect_0:SD_DAT_s1_writedata -> SD_DAT:writedata
	wire  [31:0] mm_interconnect_0_switch_pio_s1_readdata;                           // switch_pio:readdata -> mm_interconnect_0:switch_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_switch_pio_s1_address;                            // mm_interconnect_0:switch_pio_s1_address -> switch_pio:address
	wire         mm_interconnect_0_button_pio_s1_chipselect;                         // mm_interconnect_0:button_pio_s1_chipselect -> button_pio:chipselect
	wire  [31:0] mm_interconnect_0_button_pio_s1_readdata;                           // button_pio:readdata -> mm_interconnect_0:button_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_button_pio_s1_address;                            // mm_interconnect_0:button_pio_s1_address -> button_pio:address
	wire         mm_interconnect_0_button_pio_s1_write;                              // mm_interconnect_0:button_pio_s1_write -> button_pio:write_n
	wire  [31:0] mm_interconnect_0_button_pio_s1_writedata;                          // mm_interconnect_0:button_pio_s1_writedata -> button_pio:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                            // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                              // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                               // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                                 // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                             // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                            // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                              // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                               // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                 // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                             // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_uart_0_s1_chipselect;                             // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                               // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                                // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                                   // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                          // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                                  // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                              // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         mm_interconnect_0_sdram_0_s1_chipselect;                            // mm_interconnect_0:sdram_0_s1_chipselect -> sdram_0:az_cs
	wire  [15:0] mm_interconnect_0_sdram_0_s1_readdata;                              // sdram_0:za_data -> mm_interconnect_0:sdram_0_s1_readdata
	wire         mm_interconnect_0_sdram_0_s1_waitrequest;                           // sdram_0:za_waitrequest -> mm_interconnect_0:sdram_0_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_0_s1_address;                               // mm_interconnect_0:sdram_0_s1_address -> sdram_0:az_addr
	wire         mm_interconnect_0_sdram_0_s1_read;                                  // mm_interconnect_0:sdram_0_s1_read -> sdram_0:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_0_s1_byteenable;                            // mm_interconnect_0:sdram_0_s1_byteenable -> sdram_0:az_be_n
	wire         mm_interconnect_0_sdram_0_s1_readdatavalid;                         // sdram_0:za_valid -> mm_interconnect_0:sdram_0_s1_readdatavalid
	wire         mm_interconnect_0_sdram_0_s1_write;                                 // mm_interconnect_0:sdram_0_s1_write -> sdram_0:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_0_s1_writedata;                             // mm_interconnect_0:sdram_0_s1_writedata -> sdram_0:az_data
	wire   [7:0] mm_interconnect_0_cfi_flash_0_uas_readdata;                         // cfi_flash_0:uas_readdata -> mm_interconnect_0:cfi_flash_0_uas_readdata
	wire         mm_interconnect_0_cfi_flash_0_uas_waitrequest;                      // cfi_flash_0:uas_waitrequest -> mm_interconnect_0:cfi_flash_0_uas_waitrequest
	wire         mm_interconnect_0_cfi_flash_0_uas_debugaccess;                      // mm_interconnect_0:cfi_flash_0_uas_debugaccess -> cfi_flash_0:uas_debugaccess
	wire  [21:0] mm_interconnect_0_cfi_flash_0_uas_address;                          // mm_interconnect_0:cfi_flash_0_uas_address -> cfi_flash_0:uas_address
	wire         mm_interconnect_0_cfi_flash_0_uas_read;                             // mm_interconnect_0:cfi_flash_0_uas_read -> cfi_flash_0:uas_read
	wire   [0:0] mm_interconnect_0_cfi_flash_0_uas_byteenable;                       // mm_interconnect_0:cfi_flash_0_uas_byteenable -> cfi_flash_0:uas_byteenable
	wire         mm_interconnect_0_cfi_flash_0_uas_readdatavalid;                    // cfi_flash_0:uas_readdatavalid -> mm_interconnect_0:cfi_flash_0_uas_readdatavalid
	wire         mm_interconnect_0_cfi_flash_0_uas_lock;                             // mm_interconnect_0:cfi_flash_0_uas_lock -> cfi_flash_0:uas_lock
	wire         mm_interconnect_0_cfi_flash_0_uas_write;                            // mm_interconnect_0:cfi_flash_0_uas_write -> cfi_flash_0:uas_write
	wire   [7:0] mm_interconnect_0_cfi_flash_0_uas_writedata;                        // mm_interconnect_0:cfi_flash_0_uas_writedata -> cfi_flash_0:uas_writedata
	wire   [0:0] mm_interconnect_0_cfi_flash_0_uas_burstcount;                       // mm_interconnect_0:cfi_flash_0_uas_burstcount -> cfi_flash_0:uas_burstcount
	wire         irq_mapper_receiver0_irq;                                           // epcs_controller:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                           // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                           // uart_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                           // timer_0:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                           // button_pio:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                           // timer_1:irq -> irq_mapper:receiver5_irq
	wire  [31:0] nios2_qsys_0_irq_irq;                                               // irq_mapper:sender_irq -> nios2_qsys_0:irq
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [Audio_0:iRST_N, SD_CLK:reset_n, SD_CMD:reset_n, SD_DAT:reset_n, SEG7_Display:iRST_N, button_pio:reset_n, cfi_flash_0:reset_reset, epcs_controller:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, led_green:reset_n, led_red:reset_n, mm_interconnect_0:nios2_qsys_0_reset_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, rst_translator:in_reset, sdram_0:reset_n, sram_16bit_512k_0:iRST_N, switch_pio:reset_n, timer_0:reset_n, timer_1:reset_n, tri_state_bridge_0_bridge_0:reset, tri_state_bridge_0_pinSharer_0:reset_reset, uart_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                                 // rst_controller:reset_req -> [epcs_controller:reset_req, nios2_qsys_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_debug_reset_request_reset;                             // nios2_qsys_0:debug_reset_request -> rst_controller:reset_in1

	AUDIO_DAC_FIFO #(
		.REF_CLK     (18432000),
		.SAMPLE_RATE (48000),
		.DATA_WIDTH  (16),
		.CHANNEL_NUM (2)
	) audio_0 (
		.iWR_CLK   (clk_clk_in_clk),                                     //                   clk.clk
		.oAUD_DATA (audio_0_avalon_slave_0_export_oAUD_DATA),            // avalon_slave_0_export.export
		.oAUD_LRCK (audio_0_avalon_slave_0_export_oAUD_LRCK),            //                      .export
		.oAUD_BCK  (audio_0_avalon_slave_0_export_oAUD_BCK),             //                      .export
		.oAUD_XCK  (audio_0_avalon_slave_0_export_oAUD_XCK),             //                      .export
		.iCLK_18_4 (audio_0_avalon_slave_0_export_iCLK_18_4),            //                      .export
		.iDATA     (mm_interconnect_0_audio_0_avalon_slave_0_writedata), //        avalon_slave_0.writedata
		.iWR       (mm_interconnect_0_audio_0_avalon_slave_0_write),     //                      .write
		.oDATA     (mm_interconnect_0_audio_0_avalon_slave_0_readdata),  //                      .readdata
		.iRST_N    (~rst_controller_reset_out_reset)                     //               reset_n.reset_n
	);

	system_0_SD_CLK sd_clk (
		.clk        (clk_clk_in_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_sd_clk_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sd_clk_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sd_clk_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sd_clk_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sd_clk_s1_readdata),   //                    .readdata
		.out_port   (sd_clk_external_connection_export)       // external_connection.export
	);

	system_0_SD_CMD sd_cmd (
		.clk        (clk_clk_in_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_sd_cmd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sd_cmd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sd_cmd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sd_cmd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sd_cmd_s1_readdata),   //                    .readdata
		.bidir_port (sd_cmd_external_connection_export)       // external_connection.export
	);

	system_0_SD_CMD sd_dat (
		.clk        (clk_clk_in_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_sd_dat_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sd_dat_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sd_dat_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sd_dat_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sd_dat_s1_readdata),   //                    .readdata
		.bidir_port (sd_dat_external_connection_export)       // external_connection.export
	);

	SEG7_LUT_8 seg7_display (
		.iCLK   (clk_clk_in_clk),                                        //          clk.clk
		.iWR    (mm_interconnect_0_seg7_display_avalon_slave_write),     // avalon_slave.write
		.iDIG   (mm_interconnect_0_seg7_display_avalon_slave_writedata), //             .writedata
		.oSEG0  (seg7_display_conduit_end_oSEG0),                        //  conduit_end.export
		.oSEG1  (seg7_display_conduit_end_oSEG1),                        //             .export
		.oSEG2  (seg7_display_conduit_end_oSEG2),                        //             .export
		.oSEG3  (seg7_display_conduit_end_oSEG3),                        //             .export
		.oSEG4  (seg7_display_conduit_end_oSEG4),                        //             .export
		.oSEG5  (seg7_display_conduit_end_oSEG5),                        //             .export
		.oSEG6  (seg7_display_conduit_end_oSEG6),                        //             .export
		.oSEG7  (seg7_display_conduit_end_oSEG7),                        //             .export
		.iRST_N (~rst_controller_reset_out_reset)                        //      reset_n.reset_n
	);

	system_0_button_pio button_pio (
		.clk        (clk_clk_in_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_button_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_pio_s1_readdata),   //                    .readdata
		.in_port    (button_pio_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                    //                 irq.irq
	);

	system_0_cfi_flash_0 #(
		.TCM_ADDRESS_W                  (22),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (160),
		.TCM_WRITE_WAIT                 (160),
		.TCM_SETUP_WAIT                 (40),
		.TCM_DATA_HOLD                  (40),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) cfi_flash_0 (
		.clk_clk              (clk_clk_in_clk),                                  //   clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                  // reset.reset
		.uas_address          (mm_interconnect_0_cfi_flash_0_uas_address),       //   uas.address
		.uas_burstcount       (mm_interconnect_0_cfi_flash_0_uas_burstcount),    //      .burstcount
		.uas_read             (mm_interconnect_0_cfi_flash_0_uas_read),          //      .read
		.uas_write            (mm_interconnect_0_cfi_flash_0_uas_write),         //      .write
		.uas_waitrequest      (mm_interconnect_0_cfi_flash_0_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (mm_interconnect_0_cfi_flash_0_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable       (mm_interconnect_0_cfi_flash_0_uas_byteenable),    //      .byteenable
		.uas_readdata         (mm_interconnect_0_cfi_flash_0_uas_readdata),      //      .readdata
		.uas_writedata        (mm_interconnect_0_cfi_flash_0_uas_writedata),     //      .writedata
		.uas_lock             (mm_interconnect_0_cfi_flash_0_uas_lock),          //      .lock
		.uas_debugaccess      (mm_interconnect_0_cfi_flash_0_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (cfi_flash_0_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_read_n_out       (cfi_flash_0_tcm_read_n_out),                      //      .read_n_out
		.tcm_chipselect_n_out (cfi_flash_0_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_request          (cfi_flash_0_tcm_request),                         //      .request
		.tcm_grant            (cfi_flash_0_tcm_grant),                           //      .grant
		.tcm_address_out      (cfi_flash_0_tcm_address_out),                     //      .address_out
		.tcm_data_out         (cfi_flash_0_tcm_data_out),                        //      .data_out
		.tcm_data_outen       (cfi_flash_0_tcm_data_outen),                      //      .data_outen
		.tcm_data_in          (cfi_flash_0_tcm_data_in)                          //      .data_in
	);

	system_0_epcs_controller epcs_controller (
		.clk        (clk_clk_in_clk),                                                 //               clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                                //             reset.reset_n
		.reset_req  (rst_controller_reset_out_reset_req),                             //                  .reset_req
		.address    (mm_interconnect_0_epcs_controller_epcs_control_port_address),    // epcs_control_port.address
		.chipselect (mm_interconnect_0_epcs_controller_epcs_control_port_chipselect), //                  .chipselect
		.read_n     (~mm_interconnect_0_epcs_controller_epcs_control_port_read),      //                  .read_n
		.readdata   (mm_interconnect_0_epcs_controller_epcs_control_port_readdata),   //                  .readdata
		.write_n    (~mm_interconnect_0_epcs_controller_epcs_control_port_write),     //                  .write_n
		.writedata  (mm_interconnect_0_epcs_controller_epcs_control_port_writedata),  //                  .writedata
		.irq        (irq_mapper_receiver0_irq)                                        //               irq.irq
	);

	system_0_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk_in_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	system_0_led_green led_green (
		.clk        (clk_clk_in_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_led_green_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_green_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_green_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_green_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_green_s1_readdata),   //                    .readdata
		.out_port   (led_green_external_connection_export)       // external_connection.export
	);

	system_0_led_red led_red (
		.clk        (clk_clk_in_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_led_red_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_red_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_red_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_red_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_red_s1_readdata),   //                    .readdata
		.out_port   (led_red_external_connection_export)       // external_connection.export
	);

	system_0_nios2_qsys_0 nios2_qsys_0 (
		.clk                                 (clk_clk_in_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_qsys_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_qsys_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_qsys_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_qsys_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_qsys_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_qsys_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_qsys_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_qsys_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_qsys_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_qsys_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_qsys_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_qsys_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_qsys_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_qsys_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_qsys_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	system_0_sdram_0 sdram_0 (
		.clk            (clk_clk_in_clk),                             //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),            // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_0_wire_addr),                          //  wire.export
		.zs_ba          (sdram_0_wire_ba),                            //      .export
		.zs_cas_n       (sdram_0_wire_cas_n),                         //      .export
		.zs_cke         (sdram_0_wire_cke),                           //      .export
		.zs_cs_n        (sdram_0_wire_cs_n),                          //      .export
		.zs_dq          (sdram_0_wire_dq),                            //      .export
		.zs_dqm         (sdram_0_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_0_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_0_wire_we_n)                           //      .export
	);

	SRAM_16Bit_512K sram_16bit_512k_0 (
		.iCLK      (clk_clk_in_clk),                                                 //                   clk.clk
		.SRAM_DQ   (sram_16bit_512k_0_avalon_slave_0_export_DQ),                     // avalon_slave_0_export.export
		.SRAM_ADDR (sram_16bit_512k_0_avalon_slave_0_export_ADDR),                   //                      .export
		.SRAM_UB_N (sram_16bit_512k_0_avalon_slave_0_export_UB_N),                   //                      .export
		.SRAM_LB_N (sram_16bit_512k_0_avalon_slave_0_export_LB_N),                   //                      .export
		.SRAM_WE_N (sram_16bit_512k_0_avalon_slave_0_export_WE_N),                   //                      .export
		.SRAM_CE_N (sram_16bit_512k_0_avalon_slave_0_export_CE_N),                   //                      .export
		.SRAM_OE_N (sram_16bit_512k_0_avalon_slave_0_export_OE_N),                   //                      .export
		.iDATA     (mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_writedata),   //        avalon_slave_0.writedata
		.oDATA     (mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_readdata),    //                      .readdata
		.iADDR     (mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_address),     //                      .address
		.iWE_N     (~mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_write),      //                      .write_n
		.iOE_N     (~mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_read),       //                      .read_n
		.iCE_N     (~mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_chipselect), //                      .chipselect_n
		.iBE_N     (~mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_byteenable), //                      .byteenable_n
		.iRST_N    (~rst_controller_reset_out_reset)                                 //               reset_n.reset_n
	);

	system_0_switch_pio switch_pio (
		.clk      (clk_clk_in_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_switch_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switch_pio_s1_readdata), //                    .readdata
		.in_port  (switch_pio_external_connection_export)     // external_connection.export
	);

	system_0_timer_0 timer_0 (
		.clk        (clk_clk_in_clk),                          //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	system_0_timer_0 timer_1 (
		.clk        (clk_clk_in_clk),                          //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                 //   irq.irq
	);

	system_0_tri_state_bridge_0_bridge_0 tri_state_bridge_0_bridge_0 (
		.clk                               (clk_clk_in_clk),                                                     //   clk.clk
		.reset                             (rst_controller_reset_out_reset),                                     // reset.reset
		.request                           (tri_state_bridge_0_pinsharer_0_tcm_request),                         //   tcs.request
		.grant                             (tri_state_bridge_0_pinsharer_0_tcm_grant),                           //      .grant
		.tcs_tri_state_bridge_0_data       (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out),     //      .tri_state_bridge_0_data_out
		.tcs_tri_state_bridge_0_data_outen (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen),   //      .tri_state_bridge_0_data_outen
		.tcs_tri_state_bridge_0_data_in    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in),      //      .tri_state_bridge_0_data_in
		.tcs_write_n_to_the_cfi_flash_0    (tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out),  //      .write_n_to_the_cfi_flash_0_out
		.tcs_tri_state_bridge_0_readn      (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out),    //      .tri_state_bridge_0_readn_out
		.tcs_tri_state_bridge_0_address    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out),  //      .tri_state_bridge_0_address_out
		.tcs_select_n_to_the_cfi_flash_0   (tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out), //      .select_n_to_the_cfi_flash_0_out
		.tri_state_bridge_0_data           (tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_data),            //   out.tri_state_bridge_0_data
		.write_n_to_the_cfi_flash_0        (tri_state_bridge_0_bridge_0_out_write_n_to_the_cfi_flash_0),         //      .write_n_to_the_cfi_flash_0
		.tri_state_bridge_0_readn          (tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_readn),           //      .tri_state_bridge_0_readn
		.tri_state_bridge_0_address        (tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_address),         //      .tri_state_bridge_0_address
		.select_n_to_the_cfi_flash_0       (tri_state_bridge_0_bridge_0_out_select_n_to_the_cfi_flash_0)         //      .select_n_to_the_cfi_flash_0
	);

	system_0_tri_state_bridge_0_pinSharer_0 tri_state_bridge_0_pinsharer_0 (
		.clk_clk                       (clk_clk_in_clk),                                                     //   clk.clk
		.reset_reset                   (rst_controller_reset_out_reset),                                     // reset.reset
		.request                       (tri_state_bridge_0_pinsharer_0_tcm_request),                         //   tcm.request
		.grant                         (tri_state_bridge_0_pinsharer_0_tcm_grant),                           //      .grant
		.tri_state_bridge_0_address    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out),  //      .tri_state_bridge_0_address_out
		.tri_state_bridge_0_readn      (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out),    //      .tri_state_bridge_0_readn_out
		.write_n_to_the_cfi_flash_0    (tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out),  //      .write_n_to_the_cfi_flash_0_out
		.tri_state_bridge_0_data       (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out),     //      .tri_state_bridge_0_data_out
		.tri_state_bridge_0_data_in    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in),      //      .tri_state_bridge_0_data_in
		.tri_state_bridge_0_data_outen (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen),   //      .tri_state_bridge_0_data_outen
		.select_n_to_the_cfi_flash_0   (tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out), //      .select_n_to_the_cfi_flash_0_out
		.tcs0_request                  (cfi_flash_0_tcm_request),                                            //  tcs0.request
		.tcs0_grant                    (cfi_flash_0_tcm_grant),                                              //      .grant
		.tcs0_address_out              (cfi_flash_0_tcm_address_out),                                        //      .address_out
		.tcs0_read_n_out               (cfi_flash_0_tcm_read_n_out),                                         //      .read_n_out
		.tcs0_write_n_out              (cfi_flash_0_tcm_write_n_out),                                        //      .write_n_out
		.tcs0_data_out                 (cfi_flash_0_tcm_data_out),                                           //      .data_out
		.tcs0_data_in                  (cfi_flash_0_tcm_data_in),                                            //      .data_in
		.tcs0_data_outen               (cfi_flash_0_tcm_data_outen),                                         //      .data_outen
		.tcs0_chipselect_n_out         (cfi_flash_0_tcm_chipselect_n_out)                                    //      .chipselect_n_out
	);

	system_0_uart_0 uart_0 (
		.clk           (clk_clk_in_clk),                            //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (uart_0_external_connection_rxd),            // external_connection.export
		.txd           (uart_0_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver2_irq)                   //                 irq.irq
	);

	system_0_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                    (clk_clk_in_clk),                                                 //                                  clk_clk.clk
		.nios2_qsys_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                 // nios2_qsys_0_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address               (nios2_qsys_0_data_master_address),                               //                 nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest           (nios2_qsys_0_data_master_waitrequest),                           //                                         .waitrequest
		.nios2_qsys_0_data_master_byteenable            (nios2_qsys_0_data_master_byteenable),                            //                                         .byteenable
		.nios2_qsys_0_data_master_read                  (nios2_qsys_0_data_master_read),                                  //                                         .read
		.nios2_qsys_0_data_master_readdata              (nios2_qsys_0_data_master_readdata),                              //                                         .readdata
		.nios2_qsys_0_data_master_readdatavalid         (nios2_qsys_0_data_master_readdatavalid),                         //                                         .readdatavalid
		.nios2_qsys_0_data_master_write                 (nios2_qsys_0_data_master_write),                                 //                                         .write
		.nios2_qsys_0_data_master_writedata             (nios2_qsys_0_data_master_writedata),                             //                                         .writedata
		.nios2_qsys_0_data_master_debugaccess           (nios2_qsys_0_data_master_debugaccess),                           //                                         .debugaccess
		.nios2_qsys_0_instruction_master_address        (nios2_qsys_0_instruction_master_address),                        //          nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest    (nios2_qsys_0_instruction_master_waitrequest),                    //                                         .waitrequest
		.nios2_qsys_0_instruction_master_read           (nios2_qsys_0_instruction_master_read),                           //                                         .read
		.nios2_qsys_0_instruction_master_readdata       (nios2_qsys_0_instruction_master_readdata),                       //                                         .readdata
		.nios2_qsys_0_instruction_master_readdatavalid  (nios2_qsys_0_instruction_master_readdatavalid),                  //                                         .readdatavalid
		.Audio_0_avalon_slave_0_write                   (mm_interconnect_0_audio_0_avalon_slave_0_write),                 //                   Audio_0_avalon_slave_0.write
		.Audio_0_avalon_slave_0_readdata                (mm_interconnect_0_audio_0_avalon_slave_0_readdata),              //                                         .readdata
		.Audio_0_avalon_slave_0_writedata               (mm_interconnect_0_audio_0_avalon_slave_0_writedata),             //                                         .writedata
		.button_pio_s1_address                          (mm_interconnect_0_button_pio_s1_address),                        //                            button_pio_s1.address
		.button_pio_s1_write                            (mm_interconnect_0_button_pio_s1_write),                          //                                         .write
		.button_pio_s1_readdata                         (mm_interconnect_0_button_pio_s1_readdata),                       //                                         .readdata
		.button_pio_s1_writedata                        (mm_interconnect_0_button_pio_s1_writedata),                      //                                         .writedata
		.button_pio_s1_chipselect                       (mm_interconnect_0_button_pio_s1_chipselect),                     //                                         .chipselect
		.cfi_flash_0_uas_address                        (mm_interconnect_0_cfi_flash_0_uas_address),                      //                          cfi_flash_0_uas.address
		.cfi_flash_0_uas_write                          (mm_interconnect_0_cfi_flash_0_uas_write),                        //                                         .write
		.cfi_flash_0_uas_read                           (mm_interconnect_0_cfi_flash_0_uas_read),                         //                                         .read
		.cfi_flash_0_uas_readdata                       (mm_interconnect_0_cfi_flash_0_uas_readdata),                     //                                         .readdata
		.cfi_flash_0_uas_writedata                      (mm_interconnect_0_cfi_flash_0_uas_writedata),                    //                                         .writedata
		.cfi_flash_0_uas_burstcount                     (mm_interconnect_0_cfi_flash_0_uas_burstcount),                   //                                         .burstcount
		.cfi_flash_0_uas_byteenable                     (mm_interconnect_0_cfi_flash_0_uas_byteenable),                   //                                         .byteenable
		.cfi_flash_0_uas_readdatavalid                  (mm_interconnect_0_cfi_flash_0_uas_readdatavalid),                //                                         .readdatavalid
		.cfi_flash_0_uas_waitrequest                    (mm_interconnect_0_cfi_flash_0_uas_waitrequest),                  //                                         .waitrequest
		.cfi_flash_0_uas_lock                           (mm_interconnect_0_cfi_flash_0_uas_lock),                         //                                         .lock
		.cfi_flash_0_uas_debugaccess                    (mm_interconnect_0_cfi_flash_0_uas_debugaccess),                  //                                         .debugaccess
		.epcs_controller_epcs_control_port_address      (mm_interconnect_0_epcs_controller_epcs_control_port_address),    //        epcs_controller_epcs_control_port.address
		.epcs_controller_epcs_control_port_write        (mm_interconnect_0_epcs_controller_epcs_control_port_write),      //                                         .write
		.epcs_controller_epcs_control_port_read         (mm_interconnect_0_epcs_controller_epcs_control_port_read),       //                                         .read
		.epcs_controller_epcs_control_port_readdata     (mm_interconnect_0_epcs_controller_epcs_control_port_readdata),   //                                         .readdata
		.epcs_controller_epcs_control_port_writedata    (mm_interconnect_0_epcs_controller_epcs_control_port_writedata),  //                                         .writedata
		.epcs_controller_epcs_control_port_chipselect   (mm_interconnect_0_epcs_controller_epcs_control_port_chipselect), //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),        //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),          //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),           //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),       //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),      //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),    //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),     //                                         .chipselect
		.led_green_s1_address                           (mm_interconnect_0_led_green_s1_address),                         //                             led_green_s1.address
		.led_green_s1_write                             (mm_interconnect_0_led_green_s1_write),                           //                                         .write
		.led_green_s1_readdata                          (mm_interconnect_0_led_green_s1_readdata),                        //                                         .readdata
		.led_green_s1_writedata                         (mm_interconnect_0_led_green_s1_writedata),                       //                                         .writedata
		.led_green_s1_chipselect                        (mm_interconnect_0_led_green_s1_chipselect),                      //                                         .chipselect
		.led_red_s1_address                             (mm_interconnect_0_led_red_s1_address),                           //                               led_red_s1.address
		.led_red_s1_write                               (mm_interconnect_0_led_red_s1_write),                             //                                         .write
		.led_red_s1_readdata                            (mm_interconnect_0_led_red_s1_readdata),                          //                                         .readdata
		.led_red_s1_writedata                           (mm_interconnect_0_led_red_s1_writedata),                         //                                         .writedata
		.led_red_s1_chipselect                          (mm_interconnect_0_led_red_s1_chipselect),                        //                                         .chipselect
		.nios2_qsys_0_debug_mem_slave_address           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),         //             nios2_qsys_0_debug_mem_slave.address
		.nios2_qsys_0_debug_mem_slave_write             (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),           //                                         .write
		.nios2_qsys_0_debug_mem_slave_read              (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),            //                                         .read
		.nios2_qsys_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),        //                                         .readdata
		.nios2_qsys_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),       //                                         .writedata
		.nios2_qsys_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),      //                                         .byteenable
		.nios2_qsys_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest),     //                                         .waitrequest
		.nios2_qsys_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess),     //                                         .debugaccess
		.SD_CLK_s1_address                              (mm_interconnect_0_sd_clk_s1_address),                            //                                SD_CLK_s1.address
		.SD_CLK_s1_write                                (mm_interconnect_0_sd_clk_s1_write),                              //                                         .write
		.SD_CLK_s1_readdata                             (mm_interconnect_0_sd_clk_s1_readdata),                           //                                         .readdata
		.SD_CLK_s1_writedata                            (mm_interconnect_0_sd_clk_s1_writedata),                          //                                         .writedata
		.SD_CLK_s1_chipselect                           (mm_interconnect_0_sd_clk_s1_chipselect),                         //                                         .chipselect
		.SD_CMD_s1_address                              (mm_interconnect_0_sd_cmd_s1_address),                            //                                SD_CMD_s1.address
		.SD_CMD_s1_write                                (mm_interconnect_0_sd_cmd_s1_write),                              //                                         .write
		.SD_CMD_s1_readdata                             (mm_interconnect_0_sd_cmd_s1_readdata),                           //                                         .readdata
		.SD_CMD_s1_writedata                            (mm_interconnect_0_sd_cmd_s1_writedata),                          //                                         .writedata
		.SD_CMD_s1_chipselect                           (mm_interconnect_0_sd_cmd_s1_chipselect),                         //                                         .chipselect
		.SD_DAT_s1_address                              (mm_interconnect_0_sd_dat_s1_address),                            //                                SD_DAT_s1.address
		.SD_DAT_s1_write                                (mm_interconnect_0_sd_dat_s1_write),                              //                                         .write
		.SD_DAT_s1_readdata                             (mm_interconnect_0_sd_dat_s1_readdata),                           //                                         .readdata
		.SD_DAT_s1_writedata                            (mm_interconnect_0_sd_dat_s1_writedata),                          //                                         .writedata
		.SD_DAT_s1_chipselect                           (mm_interconnect_0_sd_dat_s1_chipselect),                         //                                         .chipselect
		.sdram_0_s1_address                             (mm_interconnect_0_sdram_0_s1_address),                           //                               sdram_0_s1.address
		.sdram_0_s1_write                               (mm_interconnect_0_sdram_0_s1_write),                             //                                         .write
		.sdram_0_s1_read                                (mm_interconnect_0_sdram_0_s1_read),                              //                                         .read
		.sdram_0_s1_readdata                            (mm_interconnect_0_sdram_0_s1_readdata),                          //                                         .readdata
		.sdram_0_s1_writedata                           (mm_interconnect_0_sdram_0_s1_writedata),                         //                                         .writedata
		.sdram_0_s1_byteenable                          (mm_interconnect_0_sdram_0_s1_byteenable),                        //                                         .byteenable
		.sdram_0_s1_readdatavalid                       (mm_interconnect_0_sdram_0_s1_readdatavalid),                     //                                         .readdatavalid
		.sdram_0_s1_waitrequest                         (mm_interconnect_0_sdram_0_s1_waitrequest),                       //                                         .waitrequest
		.sdram_0_s1_chipselect                          (mm_interconnect_0_sdram_0_s1_chipselect),                        //                                         .chipselect
		.SEG7_Display_avalon_slave_write                (mm_interconnect_0_seg7_display_avalon_slave_write),              //                SEG7_Display_avalon_slave.write
		.SEG7_Display_avalon_slave_writedata            (mm_interconnect_0_seg7_display_avalon_slave_writedata),          //                                         .writedata
		.sram_16bit_512k_0_avalon_slave_0_address       (mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_address),     //         sram_16bit_512k_0_avalon_slave_0.address
		.sram_16bit_512k_0_avalon_slave_0_write         (mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_write),       //                                         .write
		.sram_16bit_512k_0_avalon_slave_0_read          (mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_read),        //                                         .read
		.sram_16bit_512k_0_avalon_slave_0_readdata      (mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_readdata),    //                                         .readdata
		.sram_16bit_512k_0_avalon_slave_0_writedata     (mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_writedata),   //                                         .writedata
		.sram_16bit_512k_0_avalon_slave_0_byteenable    (mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_byteenable),  //                                         .byteenable
		.sram_16bit_512k_0_avalon_slave_0_chipselect    (mm_interconnect_0_sram_16bit_512k_0_avalon_slave_0_chipselect),  //                                         .chipselect
		.switch_pio_s1_address                          (mm_interconnect_0_switch_pio_s1_address),                        //                            switch_pio_s1.address
		.switch_pio_s1_readdata                         (mm_interconnect_0_switch_pio_s1_readdata),                       //                                         .readdata
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                           //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                             //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                          //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                         //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect),                        //                                         .chipselect
		.timer_1_s1_address                             (mm_interconnect_0_timer_1_s1_address),                           //                               timer_1_s1.address
		.timer_1_s1_write                               (mm_interconnect_0_timer_1_s1_write),                             //                                         .write
		.timer_1_s1_readdata                            (mm_interconnect_0_timer_1_s1_readdata),                          //                                         .readdata
		.timer_1_s1_writedata                           (mm_interconnect_0_timer_1_s1_writedata),                         //                                         .writedata
		.timer_1_s1_chipselect                          (mm_interconnect_0_timer_1_s1_chipselect),                        //                                         .chipselect
		.uart_0_s1_address                              (mm_interconnect_0_uart_0_s1_address),                            //                                uart_0_s1.address
		.uart_0_s1_write                                (mm_interconnect_0_uart_0_s1_write),                              //                                         .write
		.uart_0_s1_read                                 (mm_interconnect_0_uart_0_s1_read),                               //                                         .read
		.uart_0_s1_readdata                             (mm_interconnect_0_uart_0_s1_readdata),                           //                                         .readdata
		.uart_0_s1_writedata                            (mm_interconnect_0_uart_0_s1_writedata),                          //                                         .writedata
		.uart_0_s1_begintransfer                        (mm_interconnect_0_uart_0_s1_begintransfer),                      //                                         .begintransfer
		.uart_0_s1_chipselect                           (mm_interconnect_0_uart_0_s1_chipselect)                          //                                         .chipselect
	);

	system_0_irq_mapper irq_mapper (
		.clk           (clk_clk_in_clk),                 //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (nios2_qsys_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~clk_clk_in_reset_reset_n),              // reset_in0.reset
		.reset_in1      (nios2_qsys_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk_in_clk),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
